module alu #(
	parameter MSB = 7 
)(
	output signed [MSB:0] z, 
	input sel_inv_z, 
	input sel_rbo_z, 
	input sel_shl_z, 
	input sel_add, 
	input sel_inv_x, sel_inv_y, 
	input sel_zero_x, sel_zero_y, 
	input signed [MSB:0] x, y 
);

wire signed [MSB:0] x1 = sel_zero_x ? {(MSB+1){1'b0}} : x;
wire signed [MSB:0] y1 = sel_zero_y ? {(MSB+1){1'b0}} : y;
wire signed [MSB:0] x2 = sel_inv_x ? ~x1 : x1;
wire signed [MSB:0] y2 = sel_inv_y ? ~y1 : y1;
wire signed [MSB:0] z1 = sel_add ? (x2 + y2) : (x2 & y2);
wire signed [MSB:0] z2 = sel_shl_z ? z1 << 1 : z1;
wire signed [MSB:0] z2_r;
genvar i;
generate
	for(i=0;i<=MSB;i=i+1) begin :rbo_i
		assign z2_r[i] = z2[MSB-i];
	end
endgenerate
wire signed [MSB:0] z3 = sel_rbo_z ? z2_r : z2;
wire signed [MSB:0] z4 = sel_inv_z ? ~z3 : z3;
assign z = z4;

endmodule


/*
`timescale 1ps/1ps

module alu_tb;

	parameter MSB = 7 ;
	wire signed [MSB:0] z;
	reg [7:0] f;
	reg signed [MSB:0] x, y;

alu #(
	. MSB (MSB)
) u_alu(
	.z(z), 
	.sel_inv_z(f[7]), 
	.sel_rbo_z(f[6]), 
	.sel_shl_z(f[5]), 
	.sel_add(f[4]), 
	.sel_inv_x(f[3]), .sel_inv_y(f[2]), 
	.sel_zero_x(f[1]), .sel_zero_y(f[0]), 
	.x(x), .y(y) 
);

initial begin
	$dumpfile("a.fst");
	$dumpvars(0, alu_tb);
	f = 8'b00000000;
	repeat(9'b100000000) begin
		#1;
		x = $urandom_range(0, 1<<(MSB+1)-1);
		y = $urandom_range(0, 1<<(MSB+1)-1);
		f = f + 1;
	end
	$finish;
end

endmodule
*/


module cpu #(
	parameter IMSB = 15, 
	parameter PMSB = 7, 
	parameter AMSB = 7, 
	parameter DMSB = 7 
)(
	output idle, 
	input signed [DMSB:0] rdata, 
	output write, 
	output reg signed [DMSB:0] wdata, 
	output reg [AMSB:0] addr, 
	input [IMSB:0] inst, 
	output reg [PMSB:0] pc, 
	input rstn, setn, clk 
);

reg signed [DMSB:0] z;
wire signed [DMSB:0] x, y, nxt_z;
wire eq = ~|nxt_z;
wire lt = nxt_z[DMSB];
wire gt = ~|{eq,lt};

wire [1:0] src_x = inst[9:8];
assign x = 
	(src_x == 2'b11) ? wdata[DMSB:0] : 
	(src_x == 2'b01) ? addr[DMSB:0] : 
	(src_x == 2'b10) ? pc[DMSB:0] : 
	z;
wire src_y = inst[10];
assign y = 
	(src_y == 1'b1) ? rdata[DMSB:0] : 
	inst[DMSB:0];

wire ena_jmp = inst[11];
wire jeq = ena_jmp && inst[12];
wire jlt = ena_jmp && inst[13];
wire jgt = ena_jmp && inst[14];
wire jmp = |{jlt&&lt,jgt&&gt,jeq&&eq};
wire dst_pc = ena_jmp && jmp;

wire dst_wdata = ~ena_jmp && inst[12];
wire dst_addr = ~ena_jmp && inst[13];

assign write = inst[15];

assign idle = inst == 16'd0 || pc == {(PMSB+1){1'b1}};

alu #(
	. MSB (DMSB)
) u_alu(
	.z(nxt_z), 
	.sel_rbo_z(inst[7]), 
	.sel_shl_z(inst[5]), 
	.sel_inv_z(inst[5]), 
	.sel_add(inst[4]), 
	.sel_inv_x(inst[3]), .sel_inv_y(inst[2]), 
	.sel_zero_x(inst[1]), .sel_zero_y(inst[0]), 
	.x(x), .y(y) 
);

always@(negedge rstn or posedge clk) begin
	if(!rstn) z <= {(DMSB+1){1'b0}};
	else if(setn && ~idle) z <= nxt_z;
end

always@(negedge rstn or posedge clk) begin
	if(!rstn) wdata <= {(DMSB+1){1'b0}};
	else if(setn && ~idle) begin
		if(dst_wdata) wdata <= nxt_z;
	end
end

always@(negedge rstn or posedge clk) begin
	if(!rstn) addr <= {(AMSB+1){1'b0}};
	else if(setn && ~idle) begin
		if(dst_addr) addr <= nxt_z;
	end
end

always@(negedge rstn or posedge clk) begin
	if(!rstn) pc <= {(PMSB+1){1'b0}};
	else if(setn && ~idle) begin
		if(dst_pc) pc <= z;
		else pc <= pc + 1;
	end
end

endmodule


module cpu_tb_1;

reg [511:0] in_file;
reg [511:0] out_file;
integer debug_fp, in_fp, out_fp;

parameter IMSB = 15;
parameter PMSB = 7;
parameter AMSB = 7; 
parameter DMSB = 7;

reg [7:0] ram[0:(1<<AMSB)-1];
reg [AMSB:0] addr;
reg [DMSB:0] wdata, rdata;

reg [15:0] rom[0:(1<<PMSB)-1];
reg [PMSB:0] pc;
reg [IMSB:0] inst;

reg [511:0] line;
initial line = 0;
task debug_line;
	reg [PMSB:0] debug_pc;
	reg [511:0] debug_line;
	reg [7:0] debug_line_len;
	reg [7:0] debug_line_char;
	begin
		debug_fp = $fopen("a.debug","r");
		$fscanf(debug_fp, "%s\n", in_file);
		$fscanf(debug_fp, "%s\n", out_file);
		while(!$feof(debug_fp)) begin
			$fscanf(debug_fp, "%c", debug_pc);
			$fscanf(debug_fp, "%c", debug_line_len);
			debug_line = 512'd0;
			repeat(debug_line_len) begin
				$fscanf(debug_fp, "%c", debug_line_char);
				debug_line = {debug_line[511-8:0],debug_line_char};
			end
			if(pc == debug_pc) line = debug_line;
		end
		$fclose(debug_fp);
	end
endtask

reg rstn, setn, clk;

initial clk = 0;
always #1 clk = ~clk;

wire write;
wire [DMSB:0] nxt_wdata;
wire [AMSB:0] nxt_addr;
wire [PMSB:0] nxt_pc;
wire idle;

cpu #(
	.IMSB ( IMSB), 
	.PMSB ( PMSB), 
	.AMSB ( 7), 
	.DMSB ( 7 )
) u_cpu(
	.idle(idle), 
	.rdata(rdata), 
	.write(write), 
	.wdata(nxt_wdata), 
	.addr(nxt_addr), 
	.inst(inst), 
	.pc(nxt_pc), 
	.rstn(rstn), .setn(setn), .clk(clk) 
);

initial begin
	$dumpfile("a.fst");
	$dumpvars(0, cpu_tb_1);
	debug_fp = $fopen("a.debug","rb");
	$fscanf(debug_fp, "%s\n", in_file);
	$fscanf(debug_fp, "%s\n", out_file);
	$fclose(debug_fp);
	in_fp = $fopen(in_file,"r");
	out_fp = $fopen(out_file,"rb");
	rstn = 0;
	setn = 0;
	addr = 0;
	pc = 0;
	inst = 0;
	rdata = 0;
	$write("load ram\n");
	repeat(1<<(AMSB+1)) begin
		$fscanf(out_fp, "%c", wdata);
		ram[addr] = wdata;
		@(posedge clk);
		addr = addr + 1;
	end
	$write("load rom\n");
	repeat(1<<(PMSB+1)) begin
		$fscanf(out_fp, "%c", rdata);
		inst = 16'h00ff & rdata;
		$fscanf(out_fp, "%c", rdata);
		inst = (inst << 8) | (16'h00ff & rdata);
		rom[pc] = inst;
		debug_line;
		@(posedge clk);
		pc = pc + 1;
	end
	repeat(3) begin
		$write("load inst\n");
		pc = 0;
		repeat(2) @(posedge clk); rstn = 1;
		repeat(2) @(posedge clk); setn = 1;
		do begin
			addr = nxt_addr;
				wdata = nxt_wdata;
			pc = nxt_pc;
			@(posedge clk);
			if(write) rdata = ram[addr];
			inst = rom[pc];
		end while(!idle);
		repeat(2) @(posedge clk); rstn = 0;
		repeat(2) @(posedge clk); setn = 0;
	end
	$fclose(in_fp);
	$fclose(out_fp);
	$finish;
end

endmodule
